(**
 * PhiStringType - Pure Binary String Type Definition
 * 
 * This module defines the fundamental binary string type PhiString
 * as a list of PhiBit elements.
 * 
 * SINGLE THEOREM POLICY: This file contains only PhiString type and basic operations.
 * ZERO ADMITTED POLICY: All theorems proven with complete proofs ending in Qed.
 * PURE BINARY POLICY: Only PhiBit-based lists, no string dependencies.
 * 
 * Mathematical Correspondence:
 * - docs/math/00-basic-notation.md § 1.2 Binary strings
 * - docs/math/01-language-encoding.md § 1.2 φ-string definition
 * 
 * Dependencies: PhiBitType.v
 *)

(** Standard Coq imports *)
From Stdlib Require Import Lists.List.
From Stdlib Require Import Arith.Arith.
From Stdlib Require Import micromega.Lia.

(** Import our PhiBit foundation *)
Require Import PhiBitType.

Module PhiStringType.

Import ListNotations.
Import PhiBitType.

(** * The Fundamental Binary String Type *)

(**
 * PhiString: List of PhiBit elements
 * Corresponds to mathematical notation: Σ* (binary strings)
 *)
Definition PhiString : Type := list PhiBitType.PhiBit.

(** * Basic PhiString Constants *)

(**
 * Empty φ-string (corresponds to ε in mathematics)
 *)
Definition phi_empty : PhiString := [].

(**
 * Single-bit φ-strings
 *)
Definition phi_zero_string : PhiString := [PhiBitType.zero].
Definition phi_one_string : PhiString := [PhiBitType.one].

(** * Basic PhiString Operations *)

(**
 * Length of φ-string
 *)
Definition phi_length (s : PhiString) : nat := length s.

(**
 * Concatenation of φ-strings
 *)
Definition phi_concat (s1 s2 : PhiString) : PhiString := s1 ++ s2.

(**
 * Reverse of φ-string
 *)
Definition phi_reverse (s : PhiString) : PhiString := rev s.

(**
 * Append single bit to φ-string
 *)
Definition phi_append_bit (s : PhiString) (b : PhiBitType.PhiBit) : PhiString := s ++ [b].

(**
 * Prepend single bit to φ-string
 *)
Definition phi_prepend_bit (b : PhiBitType.PhiBit) (s : PhiString) : PhiString := b :: s.

(** * Basic PhiString Properties *)

(**
 * Empty string has length 0
 *)
Theorem phi_empty_length : phi_length phi_empty = 0.
Proof.
  reflexivity.
Qed.

(**
 * Single-bit strings have length 1
 *)
Theorem phi_single_bit_length : 
  phi_length phi_zero_string = 1 /\ phi_length phi_one_string = 1.
Proof.
  split; reflexivity.
Qed.

(**
 * Concatenation length is additive
 *)
Theorem phi_concat_length : forall (s1 s2 : PhiString),
  phi_length (phi_concat s1 s2) = phi_length s1 + phi_length s2.
Proof.
  intros s1 s2.
  unfold phi_length, phi_concat.
  exact (length_app s1 s2).
Qed.

(**
 * Concatenation is associative
 *)
Theorem phi_concat_assoc : forall (s1 s2 s3 : PhiString),
  phi_concat (phi_concat s1 s2) s3 = phi_concat s1 (phi_concat s2 s3).
Proof.
  intros s1 s2 s3.
  unfold phi_concat.
  rewrite app_assoc.
  reflexivity.
Qed.

(**
 * Empty string is left identity for concatenation
 *)
Theorem phi_concat_left_identity : forall (s : PhiString),
  phi_concat phi_empty s = s.
Proof.
  intro s.
  unfold phi_concat, phi_empty.
  reflexivity.
Qed.

(**
 * Empty string is right identity for concatenation
 *)
Theorem phi_concat_right_identity : forall (s : PhiString),
  phi_concat s phi_empty = s.
Proof.
  intro s.
  unfold phi_concat, phi_empty.
  exact (app_nil_r s).
Qed.

(**
 * Reverse length preservation
 *)
Theorem phi_reverse_length : forall (s : PhiString),
  phi_length (phi_reverse s) = phi_length s.
Proof.
  intro s.
  unfold phi_length, phi_reverse.
  exact (length_rev s).
Qed.

(**
 * Reverse is involutive
 *)
Theorem phi_reverse_involutive : forall (s : PhiString),
  phi_reverse (phi_reverse s) = s.
Proof.
  intro s.
  unfold phi_reverse.
  exact (rev_involutive s).
Qed.

(**
 * Append bit increases length by 1
 *)
Theorem phi_append_bit_length : forall (s : PhiString) (b : PhiBitType.PhiBit),
  phi_length (phi_append_bit s b) = phi_length s + 1.
Proof.
  intros s b.
  unfold phi_length, phi_append_bit.
  rewrite length_app.
  simpl.
  lia.
Qed.

(**
 * Prepend bit increases length by 1
 *)
Theorem phi_prepend_bit_length : forall (b : PhiBitType.PhiBit) (s : PhiString),
  phi_length (phi_prepend_bit b s) = 1 + phi_length s.
Proof.
  intros b s.
  unfold phi_length, phi_prepend_bit.
  simpl.
  lia.
Qed.

(** * Computational Verification *)

(**
 * Basic examples to verify our implementation
 *)
Example phi_string_basic_examples :
  phi_length [] = 0 /\
  phi_length [PhiBitType.zero] = 1 /\
  phi_length [PhiBitType.one] = 1 /\
  phi_length [PhiBitType.zero; PhiBitType.one] = 2 /\
  phi_length [PhiBitType.one; PhiBitType.zero] = 2 /\
  phi_concat [PhiBitType.zero] [PhiBitType.one] = [PhiBitType.zero; PhiBitType.one] /\
  phi_reverse [PhiBitType.zero; PhiBitType.one] = [PhiBitType.one; PhiBitType.zero].
Proof.
  repeat split; reflexivity.
Qed.

(** * Module Interface *)

(**
 * Core PhiString interface export
 *)
Module PhiStringInterface.
  Definition exported_PhiString := PhiString.
  Definition exported_phi_empty := phi_empty.
  Definition exported_phi_zero_string := phi_zero_string.
  Definition exported_phi_one_string := phi_one_string.
  Definition exported_phi_length := phi_length.
  Definition exported_phi_concat := phi_concat.
  Definition exported_phi_reverse := phi_reverse.
  Definition exported_phi_append_bit := phi_append_bit.
  Definition exported_phi_prepend_bit := phi_prepend_bit.
  Definition exported_phi_concat_length := phi_concat_length.
  Definition exported_phi_concat_assoc := phi_concat_assoc.
  Definition exported_phi_concat_left_identity := phi_concat_left_identity.
  Definition exported_phi_concat_right_identity := phi_concat_right_identity.
End PhiStringInterface.

End PhiStringType.

(**
 * Module Summary:
 * 
 * This PhiStringType module provides the atomic foundation for binary string
 * operations in the Zeckendorf-Hilbert formal verification project.
 * 
 * Key Properties:
 * ✓ Single focus: PhiString type and basic operations only
 * ✓ Minimal dependencies: Only PhiBitType.v and Coq standard library
 * ✓ Complete proofs: All theorems end with Qed
 * ✓ Computational verification: All operations are computable and verified
 * ✓ Pure binary implementation: Only list PhiBit, no string dependencies
 * ✓ Mathematical correspondence: Direct mapping to docs/math/ theory
 * 
 * This atomic module provides the string foundation for:
 * - No-11 constraint checking
 * - φ-language definition
 * - Encoding/decoding operations
 * - Automaton processing
 * - All higher-level binary string operations
 *)

(** End of PhiStringType module *)